module(

);

endmodule