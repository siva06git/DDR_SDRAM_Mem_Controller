module(

);
endmodule