module(
    input req_addr,
    output reg [31:0]req_write,
    output reg [31:0]req_read,
    output reg ACTIVATE,
    output reg column,
    output reg bank,
    output reg row,
    output reg req_wdata,

);

endmodule