module timing_control(
    input wire clk,
    input wire reset,

    output reg tRCD_done,
    output reg tRP_done,
    output reg tRAS_done,
    output reg tRFC_done,
    output reg tWR_done,
    output reg tWTR_done,
    output reg tRTP_done,

    

);
endmodule